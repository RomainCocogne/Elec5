package apb2wb_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "apb2wb_bridge_defines.svh"
  



endpackage