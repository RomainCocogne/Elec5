// ===============================================================================
// Copyright (c) 2015-2018 - AEDVICES Consulting
// ===============================================================================
//                     Training
//                        on
//            IP & SoC Verification Methodology
//                     using UVM
// ===============================================================================
// This material is provided as part of the training from AEDVICES Consulting,
// The directory "opencores" contains open source codes from opencores.org
// Other directories contains files and data developed by AEDVICES Consulting for
// training purposes.
// Personal copy is limited to training attendants.
// Copy and duplication other than in the context of the training is not allowed.
// ===============================================================================


// Lab : Verilog Basics - Modules and Signals
//--------------------------------------------------------------------------------
// Goals:
//  - Get started with Verilog;
//  - Be able to build a module;
//  - Be able to create a simple testbench.
//--------------------------------------------------------------------------------
// File: adder_simple.v
// Description: Module combinational addersimple, add two values and the carry in. 

module simple_adder #(parameter N = 4) (
	//LAB-TODO-STEP1-a: Define the module interface
	);

	//LAB-TODO-STEP1-b: Describe the module beharviour
endmodule