

`ifndef ADDR_WB_WIDTH
  `define ADDR_WB_WIDTH      32
`endif

`ifndef ADDR_APB_WIDTH
  `define ADDR_APB_WIDTH      32
`endif

`ifndef DATA_APB_WIDTH
  `define DATA_APB_WIDTH      32
`endif

`ifndef DATA_WB_WIDTH
  `define DATA_WB_WIDTH      32
`endif